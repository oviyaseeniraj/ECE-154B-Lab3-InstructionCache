// ucsbece154b_top_tb.v
// All Rights Reserved
// Copyright (c) 2024 UCSB ECE
// Distribution Prohibited


`define SIM

`define ASSERT(CONDITION, MESSAGE) if ((CONDITION)==1'b1); else begin $error($sformatf MESSAGE); end

module ucsbece154b_top_tb ();

// test bench contents
reg clk = 1;
always #1 clk <= ~clk;
reg reset;

integer jumptotal = 0;
integer jumppredictedcorrectly = 0;
integer branchtotal = 0;
integer branchpredictedcorrectly = 0;

// HIT/MISS TRACKING
integer total_fetches = 0;
integer icachehits = 0;
integer icachemisses = 0;
integer last_ready = 0;

ucsbece154b_top top (
    .clk(clk), .reset(reset)
);

wire [31:0] reg_zero = top.riscv.dp.rf.zero;
wire [31:0] reg_ra = top.riscv.dp.rf.ra;
wire [31:0] reg_sp = top.riscv.dp.rf.sp;
wire [31:0] reg_gp = top.riscv.dp.rf.gp;
wire [31:0] reg_tp = top.riscv.dp.rf.tp;
wire [31:0] reg_t0 = top.riscv.dp.rf.t0;
wire [31:0] reg_t1 = top.riscv.dp.rf.t1;
wire [31:0] reg_t2 = top.riscv.dp.rf.t2;
wire [31:0] reg_s0 = top.riscv.dp.rf.s0;
wire [31:0] reg_s1 = top.riscv.dp.rf.s1;
wire [31:0] reg_a0 = top.riscv.dp.rf.a0;
wire [31:0] reg_a1 = top.riscv.dp.rf.a1;
wire [31:0] reg_a2 = top.riscv.dp.rf.a2;
wire [31:0] reg_a3 = top.riscv.dp.rf.a3;
wire [31:0] reg_a4 = top.riscv.dp.rf.a4;
wire [31:0] reg_a5 = top.riscv.dp.rf.a5;
wire [31:0] reg_a6 = top.riscv.dp.rf.a6;
wire [31:0] reg_a7 = top.riscv.dp.rf.a7;
wire [31:0] reg_s2 = top.riscv.dp.rf.s2;
wire [31:0] reg_s3 = top.riscv.dp.rf.s3;
wire [31:0] reg_s4 = top.riscv.dp.rf.s4;
wire [31:0] reg_s5 = top.riscv.dp.rf.s5;
wire [31:0] reg_s6 = top.riscv.dp.rf.s6;
wire [31:0] reg_s7 = top.riscv.dp.rf.s7;
wire [31:0] reg_s8 = top.riscv.dp.rf.s8;
wire [31:0] reg_s9 = top.riscv.dp.rf.s9;
wire [31:0] reg_s10 = top.riscv.dp.rf.s10;
wire [31:0] reg_s11 = top.riscv.dp.rf.s11;
wire [31:0] reg_t3 = top.riscv.dp.rf.t3;
wire [31:0] reg_t4 = top.riscv.dp.rf.t4;
wire [31:0] reg_t5 = top.riscv.dp.rf.t5;
wire [31:0] reg_t6 = top.riscv.dp.rf.t6;

 wire [31:0] fetchpc = top.riscv.dp.PCPlus4W;

// wire [31:0] MEM_10000000 = top.dmem.DATA[6'd0];

//

integer i;
initial begin
    $display( "Begin simulation." );
    //\\ =========================== \\//

    reset = 1;
    @(negedge clk);
    @(negedge clk);
    reset = 0;
    reg prev_ready = 0;


    // Test for program 
    for (i = 0; i < 10000; i=i+1) begin
        @(negedge clk);

        if (top.icache.ReadEnable == 1 && top.icache.Ready == 1 && prev_ready == 0) begin
            total_fetches = total_fetches + 1;
            if (top.icache.MemReadRequest == 1)
                icachemisses = icachemisses + 1;
            else
                icachehits = icachehits + 1;
        end
        prev_ready = top.icache.Ready;
    // counter for jumps

        // if(top.riscv.dp.BranchE_i) branchtotal++;
        // if(top.riscv.dp.JumpE_i) jumptotal++;
        // if(~top.riscv.dp.MisspredictE_o & top.riscv.dp.BranchE_i) branchpredictedcorrectly++;
        // if(~top.riscv.dp.MisspredictE_o & top.riscv.dp.JumpE_i) jumppredictedcorrectly++;

    // counter for branches

    //         if(fetchpc==32'h00010068) begin
    //		$display("#cycles = %d", i);  
    //	 break;
    //	 end
        
    // `ASSERT(fetchpc == 32'h00010064, ("reached last instruction"));    


    // WRITE YOUR TEST HERE

    // `ASSERT(rg_zero==32'b0, ("reg_zero incorrect"));
    // `ASSERT(MEM_10000070==32'hBEEF000, ("mem.DATA[29] //incorrect"));


    //\\ =========================== \\//
        $display( "Total fetches: %d", total_fetches);
        $display( "Total icache hits: %d", icachehits);
        $display( "Total icache misses: %d", icachemisses);
        $display( "Instruction cache hit rate: %f", (icachehits*100)/total_fetches);
        $display( "Instruction cache miss rate: %f", (icachemisses*100)/total_fetches);
        $display( "End simulation.");
        $stop;
    end
end

endmodule

`undef ASSERT
